
-- 
-- Definition of  DSP48E1
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity DSP48E1 is 
   generic (ACASCREG : INTEGER := 1;
      ADREG : INTEGER := 1;
      ALUMODEREG : INTEGER := 1;
      AREG : INTEGER := 1;
      AUTORESET_PATDET : STRING := "NO_RESET";
      A_INPUT : STRING := "DIRECT";
      BCASCREG : INTEGER := 1;
      BREG : INTEGER := 1;
      B_INPUT : STRING := "DIRECT";
      CARRYINREG : INTEGER := 1;
      CARRYINSELREG : INTEGER := 1;
      CREG : INTEGER := 1;
      DREG : INTEGER := 1;
      INMODEREG : INTEGER := 1;
      IS_ALUMODE_INVERTED : BIT_VECTOR := X"0000"
      ;
      IS_CARRYIN_INVERTED : BIT := '0';
      IS_CLK_INVERTED : BIT := '0'
      ;
      IS_INMODE_INVERTED : BIT_VECTOR := X"00000"
      ;
      IS_OPMODE_INVERTED : BIT_VECTOR := X"0000000"
      ;
      MASK : BIT_VECTOR := X"3FFFFFFFFFFF";
      MREG : INTEGER := 1;
      OPMODEREG : INTEGER := 1;
      PATTERN : BIT_VECTOR := X"000000000000";
      PREG : INTEGER := 1;
      SEL_MASK : STRING := "MASK";
      SEL_PATTERN : STRING := "PATTERN";
      USE_DPORT : BOOLEAN := FALSE;
      USE_MULT : STRING := "MULTIPLY"
      ;
      USE_PATTERN_DETECT : STRING := "NO_PATDET"
      ;
      USE_SIMD : STRING := "ONE48") ;
   
   port (
      ACOUT : OUT std_logic_vector (29 DOWNTO 0) ;
      BCOUT : OUT std_logic_vector (17 DOWNTO 0) ;
      CARRYCASCOUT : OUT std_logic ;
      CARRYOUT : OUT std_logic_vector (3 DOWNTO 0) ;
      MULTSIGNOUT : OUT std_logic ;
      OVERFLOW : OUT std_logic ;
      P : OUT std_logic_vector (47 DOWNTO 0) ;
      PATTERNBDETECT : OUT std_logic ;
      PATTERNDETECT : OUT std_logic ;
      PCOUT : OUT std_logic_vector (47 DOWNTO 0) ;
      UNDERFLOW : OUT std_logic ;
      A : IN std_logic_vector (29 DOWNTO 0) ;
      ACIN : IN std_logic_vector (29 DOWNTO 0) ;
      ALUMODE : IN std_logic_vector (3 DOWNTO 0) ;
      B : IN std_logic_vector (17 DOWNTO 0) ;
      BCIN : IN std_logic_vector (17 DOWNTO 0) ;
      C : IN std_logic_vector (47 DOWNTO 0) ;
      CARRYCASCIN : IN std_logic ;
      CARRYIN : IN std_logic ;
      CARRYINSEL : IN std_logic_vector (2 DOWNTO 0) ;
      CEA1 : IN std_logic ;
      CEA2 : IN std_logic ;
      CEAD : IN std_logic ;
      CEALUMODE : IN std_logic ;
      CEB1 : IN std_logic ;
      CEB2 : IN std_logic ;
      CEC : IN std_logic ;
      CECARRYIN : IN std_logic ;
      CECTRL : IN std_logic ;
      CED : IN std_logic ;
      CEINMODE : IN std_logic ;
      CEM : IN std_logic ;
      CEP : IN std_logic ;
      CLK : IN std_logic ;
      D : IN std_logic_vector (24 DOWNTO 0) ;
      INMODE : IN std_logic_vector (4 DOWNTO 0) ;
      MULTSIGNIN : IN std_logic ;
      OPMODE : IN std_logic_vector (6 DOWNTO 0) ;
      PCIN : IN std_logic_vector (47 DOWNTO 0) ;
      RSTA : IN std_logic ;
      RSTALLCARRYIN : IN std_logic ;
      RSTALUMODE : IN std_logic ;
      RSTB : IN std_logic ;
      RSTC : IN std_logic ;
      RSTCTRL : IN std_logic ;
      RSTD : IN std_logic ;
      RSTINMODE : IN std_logic ;
      RSTM : IN std_logic ;
      RSTP : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      DSP48E1 : entity is true;
      end DSP48E1 ;

architecture NETLIST of DSP48E1 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  DSP48A1
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity DSP48A1 is 
   generic (A0REG : integer := 0;
      A1REG : integer := 1;
      B0REG : integer := 0;
      B1REG : integer := 1;
      CARRYINREG : integer := 1;
      CARRYINSEL : string := "OPMODE5";
      CARRYOUTREG : integer := 1;
      CREG : integer := 1;
      DREG : integer := 1;
      MREG : integer := 1;
      OPMODEREG : integer := 1;
      PREG : integer := 1;
      RSTTYPE : string := "SYNC") ;
   
   port (
      BCOUT : OUT std_logic_vector (17 DOWNTO 0) ;
      CARRYOUT : OUT std_logic ;
      CARRYOUTF : OUT std_logic ;
      M : OUT std_logic_vector (35 DOWNTO 0) ;
      P : OUT std_logic_vector (47 DOWNTO 0) ;
      PCOUT : OUT std_logic_vector (47 DOWNTO 0) ;
      A : IN std_logic_vector (17 DOWNTO 0) ;
      B : IN std_logic_vector (17 DOWNTO 0) ;
      C : IN std_logic_vector (47 DOWNTO 0) ;
      CARRYIN : IN std_logic ;
      CEA : IN std_logic ;
      CEB : IN std_logic ;
      CEC : IN std_logic ;
      CECARRYIN : IN std_logic ;
      CED : IN std_logic ;
      CEM : IN std_logic ;
      CEOPMODE : IN std_logic ;
      CEP : IN std_logic ;
      CLK : IN std_logic ;
      D : IN std_logic_vector (17 DOWNTO 0) ;
      OPMODE : IN std_logic_vector (7 DOWNTO 0) ;
      PCIN : IN std_logic_vector (47 DOWNTO 0) ;
      RSTA : IN std_logic ;
      RSTB : IN std_logic ;
      RSTC : IN std_logic ;
      RSTCARRYIN : IN std_logic ;
      RSTD : IN std_logic ;
      RSTM : IN std_logic ;
      RSTOPMODE : IN std_logic ;
      RSTP : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      DSP48A1 : entity is true;
      end DSP48A1 ;

architecture NETLIST of DSP48A1 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  DSP48E
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity DSP48E is 
   generic (ACASCREG : INTEGER := 1;
      ALUMODEREG : INTEGER := 1;
      AREG : INTEGER := 1;
      AUTORESET_PATTERN_DETECT : STRING := "FALSE"
      ;
      AUTORESET_PATTERN_DETECT_OPTINV : STRING := "MATCH"
      ;
      A_INPUT : STRING := "DIRECT";
      BCASCREG : INTEGER := 1;
      BREG : INTEGER := 1;
      B_INPUT : STRING := "DIRECT";
      CARRYINREG : INTEGER := 1;
      CARRYINSELREG : INTEGER := 1;
      CREG : INTEGER := 1
      ;
      MASK : BIT_VECTOR := X"001111111111111111111111111111111111111111111111"
      ;
      MREG : INTEGER := 1;
      MULTCARRYINREG : INTEGER := 1;
      OPMODEREG : INTEGER := 1
      ;
      PATTERN : BIT_VECTOR := X"000000000000000000000000000000000000000000000000"
      ;
      PREG : INTEGER := 1;
      SEL_MASK : STRING := "MASK";
      SEL_PATTERN : STRING := "PATTERN"
      ;
      SEL_ROUNDING_MASK : STRING := "SEL_MASK";
      SIM_MODE : STRING := "SAFE";
      USE_MULT : STRING := "MULT_S"
      ;
      USE_PATTERN_DETECT : STRING := "NO_PATDET"
      ;
      USE_SIMD : STRING := "ONE48") ;
   
   port (
      ACOUT : OUT std_logic_vector (29 DOWNTO 0) ;
      BCOUT : OUT std_logic_vector (17 DOWNTO 0) ;
      CARRYCASCOUT : OUT std_logic ;
      CARRYOUT : OUT std_logic_vector (3 DOWNTO 0) ;
      MULTSIGNOUT : OUT std_logic ;
      OVERFLOW : OUT std_logic ;
      P : OUT std_logic_vector (47 DOWNTO 0) ;
      PATTERNBDETECT : OUT std_logic ;
      PATTERNDETECT : OUT std_logic ;
      PCOUT : OUT std_logic_vector (47 DOWNTO 0) ;
      UNDERFLOW : OUT std_logic ;
      A : IN std_logic_vector (29 DOWNTO 0) ;
      ACIN : IN std_logic_vector (29 DOWNTO 0) ;
      ALUMODE : IN std_logic_vector (3 DOWNTO 0) ;
      B : IN std_logic_vector (17 DOWNTO 0) ;
      BCIN : IN std_logic_vector (17 DOWNTO 0) ;
      C : IN std_logic_vector (47 DOWNTO 0) ;
      CARRYCASCIN : IN std_logic ;
      CARRYIN : IN std_logic ;
      CARRYINSEL : IN std_logic_vector (2 DOWNTO 0) ;
      CEA1 : IN std_logic ;
      CEA2 : IN std_logic ;
      CEALUMODE : IN std_logic ;
      CEB1 : IN std_logic ;
      CEB2 : IN std_logic ;
      CEC : IN std_logic ;
      CECARRYIN : IN std_logic ;
      CECTRL : IN std_logic ;
      CEM : IN std_logic ;
      CEMULTCARRYIN : IN std_logic ;
      CEP : IN std_logic ;
      CLK : IN std_logic ;
      MULTSIGNIN : IN std_logic ;
      OPMODE : IN std_logic_vector (6 DOWNTO 0) ;
      PCIN : IN std_logic_vector (47 DOWNTO 0) ;
      RSTA : IN std_logic ;
      RSTALLCARRYIN : IN std_logic ;
      RSTALUMODE : IN std_logic ;
      RSTB : IN std_logic ;
      RSTC : IN std_logic ;
      RSTCTRL : IN std_logic ;
      RSTM : IN std_logic ;
      RSTP : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      DSP48E : entity is true;
      end DSP48E ;

architecture NETLIST of DSP48E is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  RAMB18
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity RAMB18 is 
   generic (DOA_REG : INTEGER := 0;
      DOB_REG : INTEGER := 0
      ;
      INITP_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_10 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_11 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_12 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_13 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_14 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_15 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_16 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_17 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_18 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_19 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_20 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_21 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_22 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_23 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_24 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_25 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_26 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_27 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_28 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_29 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_30 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_31 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_32 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_33 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_34 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_35 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_36 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_37 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_38 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_39 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_A : BIT_VECTOR := X"000000000000000000"
      ;
      INIT_B : BIT_VECTOR := X"000000000000000000"
      ;
      INIT_FILE : STRING := "NONE";
      READ_WIDTH_A : INTEGER := 0;
      READ_WIDTH_B : INTEGER := 0;
      SIM_COLLISION_CHECK : STRING := "ALL";
      SIM_MODE : STRING := "SAFE"
      ;
      SRVAL_A : BIT_VECTOR := X"000000000000000000"
      ;
      SRVAL_B : BIT_VECTOR := X"000000000000000000"
      ;
      WRITE_MODE_A : STRING := "WRITE_FIRST"
      ;
      WRITE_MODE_B : STRING := "WRITE_FIRST";
      WRITE_WIDTH_A : INTEGER := 0;
      WRITE_WIDTH_B : INTEGER := 0) ;
   
   port (
      DOA : OUT std_logic_vector (15 DOWNTO 0) ;
      DOB : OUT std_logic_vector (15 DOWNTO 0) ;
      DOPA : OUT std_logic_vector (1 DOWNTO 0) ;
      DOPB : OUT std_logic_vector (1 DOWNTO 0) ;
      ADDRA : IN std_logic_vector (13 DOWNTO 0) ;
      ADDRB : IN std_logic_vector (13 DOWNTO 0) ;
      CLKA : IN std_logic ;
      CLKB : IN std_logic ;
      DIA : IN std_logic_vector (15 DOWNTO 0) ;
      DIB : IN std_logic_vector (15 DOWNTO 0) ;
      DIPA : IN std_logic_vector (1 DOWNTO 0) ;
      DIPB : IN std_logic_vector (1 DOWNTO 0) ;
      ENA : IN std_logic ;
      ENB : IN std_logic ;
      REGCEA : IN std_logic ;
      REGCEB : IN std_logic ;
      SSRA : IN std_logic ;
      SSRB : IN std_logic ;
      WEA : IN std_logic_vector (1 DOWNTO 0) ;
      WEB : IN std_logic_vector (1 DOWNTO 0)) ;
   attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      RAMB18 : entity is true;
      end RAMB18 ;

architecture NETLIST of RAMB18 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  RAMB18SDP
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity RAMB18SDP is 
   generic (DO_REG : INTEGER := 0
      ;
      INIT : BIT_VECTOR := X"000000000000000000000000000000000000"
      ;
      INITP_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_10 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_11 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_12 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_13 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_14 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_15 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_16 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_17 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_18 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_19 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_20 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_21 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_22 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_23 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_24 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_25 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_26 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_27 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_28 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_29 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_30 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_31 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_32 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_33 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_34 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_35 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_36 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_37 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_38 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_39 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_FILE : STRING := "NONE";
      SIM_COLLISION_CHECK : STRING := "ALL";
      SIM_MODE : STRING := "SAFE"
      ;
      SRVAL : BIT_VECTOR := X"000000000000000000000000000000000000") ;
   
   port (
      DO : OUT std_logic_vector (31 DOWNTO 0) ;
      DOP : OUT std_logic_vector (3 DOWNTO 0) ;
      DI : IN std_logic_vector (31 DOWNTO 0) ;
      DIP : IN std_logic_vector (3 DOWNTO 0) ;
      RDADDR : IN std_logic_vector (8 DOWNTO 0) ;
      RDCLK : IN std_logic ;
      RDEN : IN std_logic ;
      REGCE : IN std_logic ;
      SSR : IN std_logic ;
      WE : IN std_logic_vector (3 DOWNTO 0) ;
      WRADDR : IN std_logic_vector (8 DOWNTO 0) ;
      WRCLK : IN std_logic ;
      WREN : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      RAMB18SDP : entity is true;
      end RAMB18SDP ;

architecture NETLIST of RAMB18SDP is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  RAMB36
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity RAMB36 is 
   generic (DOA_REG : integer := 0;
      DOB_REG : integer := 0
      ;
      INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_A : bit_vector := X"000000000"
      ;
      INIT_B : bit_vector := X"000000000";
      INIT_FILE : string := "NONE";
      RAM_EXTENSION_A : string := "NONE";
      RAM_EXTENSION_B : string := "NONE";
      READ_WIDTH_A : integer := 0;
      READ_WIDTH_B : integer := 0;
      SIM_COLLISION_CHECK : string := "ALL";
      SIM_MODE : string := "SAFE";
      SRVAL_A : bit_vector := X"000000000"
      ;
      SRVAL_B : bit_vector := X"000000000"
      ;
      WRITE_MODE_A : string := "WRITE_FIRST"
      ;
      WRITE_MODE_B : string := "WRITE_FIRST";
      WRITE_WIDTH_A : integer := 0;
      WRITE_WIDTH_B : integer := 0) ;
   
   port (
      CASCADEOUTLATA : OUT std_logic ;
      CASCADEOUTLATB : OUT std_logic ;
      CASCADEOUTREGA : OUT std_logic ;
      CASCADEOUTREGB : OUT std_logic ;
      DOA : OUT std_logic_vector (31 DOWNTO 0) ;
      DOB : OUT std_logic_vector (31 DOWNTO 0) ;
      DOPA : OUT std_logic_vector (3 DOWNTO 0) ;
      DOPB : OUT std_logic_vector (3 DOWNTO 0) ;
      ADDRA : IN std_logic_vector (15 DOWNTO 0) ;
      ADDRB : IN std_logic_vector (15 DOWNTO 0) ;
      CASCADEINLATA : IN std_logic ;
      CASCADEINLATB : IN std_logic ;
      CASCADEINREGA : IN std_logic ;
      CASCADEINREGB : IN std_logic ;
      CLKA : IN std_logic ;
      CLKB : IN std_logic ;
      DIA : IN std_logic_vector (31 DOWNTO 0) ;
      DIB : IN std_logic_vector (31 DOWNTO 0) ;
      DIPA : IN std_logic_vector (3 DOWNTO 0) ;
      DIPB : IN std_logic_vector (3 DOWNTO 0) ;
      ENA : IN std_logic ;
      ENB : IN std_logic ;
      REGCEA : IN std_logic ;
      REGCEB : IN std_logic ;
      SSRA : IN std_logic ;
      SSRB : IN std_logic ;
      WEA : IN std_logic_vector (3 DOWNTO 0) ;
      WEB : IN std_logic_vector (3 DOWNTO 0)) ;
   attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      RAMB36 : entity is true;
      end RAMB36 ;

architecture NETLIST of RAMB36 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  RAMB36SDP
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity RAMB36SDP is 
   generic (DO_REG : integer := 0;
      EN_ECC_READ : boolean := FALSE;
      EN_ECC_SCRUB : boolean := FALSE;
      EN_ECC_WRITE : boolean := FALSE
      ;
      INIT : bit_vector := X"000000000000000000"
      ;
      INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_FILE : string := "NONE";
      SIM_COLLISION_CHECK : string := "ALL";
      SIM_MODE : string := "SAFE"
      ;
      SRVAL : bit_vector := X"000000000000000000") ;
   
   port (
      DBITERR : OUT std_logic ;
      DO : OUT std_logic_vector (63 DOWNTO 0) ;
      DOP : OUT std_logic_vector (7 DOWNTO 0) ;
      ECCPARITY : OUT std_logic_vector (7 DOWNTO 0) ;
      SBITERR : OUT std_logic ;
      DI : IN std_logic_vector (63 DOWNTO 0) ;
      DIP : IN std_logic_vector (7 DOWNTO 0) ;
      RDADDR : IN std_logic_vector (8 DOWNTO 0) ;
      RDCLK : IN std_logic ;
      RDEN : IN std_logic ;
      REGCE : IN std_logic ;
      SSR : IN std_logic ;
      WE : IN std_logic_vector (7 DOWNTO 0) ;
      WRADDR : IN std_logic_vector (8 DOWNTO 0) ;
      WRCLK : IN std_logic ;
      WREN : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      RAMB36SDP : entity is true;
      end RAMB36SDP ;

architecture NETLIST of RAMB36SDP is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  RAMB18E1
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity RAMB18E1 is 
   generic (DOA_REG : INTEGER := 0;
      DOB_REG : INTEGER := 0
      ;
      INITP_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_10 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_11 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_12 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_13 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_14 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_15 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_16 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_17 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_18 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_19 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_20 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_21 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_22 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_23 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_24 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_25 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_26 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_27 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_28 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_29 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_30 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_31 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_32 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_33 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_34 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_35 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_36 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_37 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_38 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_39 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_A : BIT_VECTOR := X"00000";
      INIT_B : BIT_VECTOR := X"00000";
      INIT_FILE : STRING := "NONE";
      IS_CLKARDCLK_INVERTED : BIT := '0';
      IS_CLKBWRCLK_INVERTED : BIT := '0';
      IS_ENARDEN_INVERTED : BIT := '0';
      IS_ENBWREN_INVERTED : BIT := '0'
      ;
      IS_RSTRAMARSTRAM_INVERTED : BIT := '0'
      ;
      IS_RSTRAMB_INVERTED : BIT := '0'
      ;
      IS_RSTREGARSTREG_INVERTED : BIT := '0'
      ;
      IS_RSTREGB_INVERTED : BIT := '0';
      RAM_MODE : STRING := "TDP"
      ;
      RDADDR_COLLISION_HWCONFIG : STRING := "DELAYED_WRITE"
      ;
      READ_WIDTH_A : INTEGER := 0;
      READ_WIDTH_B : INTEGER := 0;
      RSTREG_PRIORITY_A : STRING := "RSTREG"
      ;
      RSTREG_PRIORITY_B : STRING := "RSTREG"
      ;
      SIM_COLLISION_CHECK : STRING := "ALL"
      ;
      SIM_DEVICE : STRING := "7SERIES";
      SRVAL_A : BIT_VECTOR := X"00000";
      SRVAL_B : BIT_VECTOR := X"00000"
      ;
      WRITE_MODE_A : STRING := "WRITE_FIRST"
      ;
      WRITE_MODE_B : STRING := "WRITE_FIRST";
      WRITE_WIDTH_A : INTEGER := 0;
      WRITE_WIDTH_B : INTEGER := 0) ;
   
   port (
      DOADO : OUT std_logic_vector (15 DOWNTO 0) ;
      DOBDO : OUT std_logic_vector (15 DOWNTO 0) ;
      DOPADOP : OUT std_logic_vector (1 DOWNTO 0) ;
      DOPBDOP : OUT std_logic_vector (1 DOWNTO 0) ;
      ADDRARDADDR : IN std_logic_vector (13 DOWNTO 0) ;
      ADDRBWRADDR : IN std_logic_vector (13 DOWNTO 0) ;
      CLKARDCLK : IN std_logic ;
      CLKBWRCLK : IN std_logic ;
      DIADI : IN std_logic_vector (15 DOWNTO 0) ;
      DIBDI : IN std_logic_vector (15 DOWNTO 0) ;
      DIPADIP : IN std_logic_vector (1 DOWNTO 0) ;
      DIPBDIP : IN std_logic_vector (1 DOWNTO 0) ;
      ENARDEN : IN std_logic ;
      ENBWREN : IN std_logic ;
      REGCEAREGCE : IN std_logic ;
      REGCEB : IN std_logic ;
      RSTRAMARSTRAM : IN std_logic ;
      RSTRAMB : IN std_logic ;
      RSTREGARSTREG : IN std_logic ;
      RSTREGB : IN std_logic ;
      WEA : IN std_logic_vector (1 DOWNTO 0) ;
      WEBWE : IN std_logic_vector (3 DOWNTO 0)) ;
   attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      RAMB18E1 : entity is true;
      end RAMB18E1 ;

architecture NETLIST of RAMB18E1 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  RAMB36E1
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity RAMB36E1 is 
   generic (DOA_REG : INTEGER := 0;
      DOB_REG : INTEGER := 0;
      EN_ECC_READ : STRING := "FALSE";
      EN_ECC_WRITE : STRING := "FALSE"
      ;
      INITP_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_10 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_11 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_12 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_13 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_14 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_15 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_16 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_17 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_18 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_19 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_20 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_21 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_22 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_23 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_24 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_25 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_26 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_27 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_28 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_29 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_30 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_31 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_32 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_33 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_34 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_35 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_36 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_37 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_38 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_39 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_40 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_41 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_42 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_43 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_44 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_45 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_46 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_47 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_48 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_49 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_4F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_50 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_51 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_52 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_53 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_54 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_55 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_56 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_57 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_58 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_59 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_5F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_60 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_61 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_62 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_63 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_64 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_65 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_66 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_67 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_68 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_69 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_6F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_70 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_71 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_72 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_73 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_74 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_75 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_76 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_77 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_78 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_79 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_7F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_A : BIT_VECTOR := X"000000000000000000000000000000000000"
      ;
      INIT_B : BIT_VECTOR := X"000000000000000000000000000000000000"
      ;
      INIT_FILE : STRING := "NONE"
      ;
      IS_CLKARDCLK_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_CLKBWRCLK_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_ENARDEN_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_ENBWREN_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_RSTRAMARSTRAM_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_RSTRAMB_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_RSTREGARSTREG_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_RSTREGB_INVERTED : BIT_VECTOR := X"0"
      ;
      RAM_EXTENSION_A : STRING := "NONE";
      RAM_EXTENSION_B : STRING := "NONE";
      RAM_MODE : STRING := "TDP"
      ;
      RDADDR_COLLISION_HWCONFIG : STRING := "DELAYED_WRITE"
      ;
      READ_WIDTH_A : INTEGER := 0;
      READ_WIDTH_B : INTEGER := 0;
      RSTREG_PRIORITY_A : STRING := "RSTREG"
      ;
      RSTREG_PRIORITY_B : STRING := "RSTREG"
      ;
      SIM_COLLISION_CHECK : STRING := "ALL"
      ;
      SIM_DEVICE : STRING := "7SERIES"
      ;
      SRVAL_A : BIT_VECTOR := X"000000000000000000000000000000000000"
      ;
      SRVAL_B : BIT_VECTOR := X"000000000000000000000000000000000000"
      ;
      WRITE_MODE_A : STRING := "WRITE_FIRST"
      ;
      WRITE_MODE_B : STRING := "WRITE_FIRST";
      WRITE_WIDTH_A : INTEGER := 0;
      WRITE_WIDTH_B : INTEGER := 0) ;
   
   port (
      CASCADEOUTA : OUT std_logic ;
      CASCADEOUTB : OUT std_logic ;
      DBITERR : OUT std_logic ;
      DOADO : OUT std_logic_vector (31 DOWNTO 0) ;
      DOBDO : OUT std_logic_vector (31 DOWNTO 0) ;
      DOPADOP : OUT std_logic_vector (3 DOWNTO 0) ;
      DOPBDOP : OUT std_logic_vector (3 DOWNTO 0) ;
      ECCPARITY : OUT std_logic_vector (7 DOWNTO 0) ;
      RDADDRECC : OUT std_logic_vector (8 DOWNTO 0) ;
      SBITERR : OUT std_logic ;
      ADDRARDADDR : IN std_logic_vector (15 DOWNTO 0) ;
      ADDRBWRADDR : IN std_logic_vector (15 DOWNTO 0) ;
      CASCADEINA : IN std_logic ;
      CASCADEINB : IN std_logic ;
      CLKARDCLK : IN std_logic ;
      CLKBWRCLK : IN std_logic ;
      DIADI : IN std_logic_vector (31 DOWNTO 0) ;
      DIBDI : IN std_logic_vector (31 DOWNTO 0) ;
      DIPADIP : IN std_logic_vector (3 DOWNTO 0) ;
      DIPBDIP : IN std_logic_vector (3 DOWNTO 0) ;
      ENARDEN : IN std_logic ;
      ENBWREN : IN std_logic ;
      INJECTDBITERR : IN std_logic ;
      INJECTSBITERR : IN std_logic ;
      REGCEAREGCE : IN std_logic ;
      REGCEB : IN std_logic ;
      RSTRAMARSTRAM : IN std_logic ;
      RSTRAMB : IN std_logic ;
      RSTREGARSTREG : IN std_logic ;
      RSTREGB : IN std_logic ;
      WEA : IN std_logic_vector (3 DOWNTO 0) ;
      WEBWE : IN std_logic_vector (7 DOWNTO 0)) ;
   attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      RAMB36E1 : entity is true;
      end RAMB36E1 ;

architecture NETLIST of RAMB36E1 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  RAMB8BWER
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity RAMB8BWER is 
   generic (DATA_WIDTH_A : integer := 0;
      DATA_WIDTH_B : integer := 0;
      DOA_REG : integer := 0;
      DOB_REG : integer := 0;
      EN_RSTRAM_A : boolean := TRUE;
      EN_RSTRAM_B : boolean := TRUE
      ;
      INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_A : bit_vector := X"00000";
      INIT_B : bit_vector := X"00000";
      INIT_FILE : string := "NONE";
      RAM_MODE : string := "TDP";
      RSTTYPE : string := "SYNC";
      RST_PRIORITY_A : string := "SR";
      RST_PRIORITY_B : string := "SR";
      SETUP_ALL : time := 1000000 ns;
      SETUP_READ_FIRST : time := 3000000 ns
      ;
      SIM_COLLISION_CHECK : string := "ALL"
      ;
      SRVAL_A : bit_vector := X"00000";
      SRVAL_B : bit_vector := X"00000"
      ;
      WRITE_MODE_A : string := "WRITE_FIRST"
      ;
      WRITE_MODE_B : string := "WRITE_FIRST") ;
   
   port (
      DOADO : OUT std_logic_vector (15 DOWNTO 0) ;
      DOBDO : OUT std_logic_vector (15 DOWNTO 0) ;
      DOPADOP : OUT std_logic_vector (1 DOWNTO 0) ;
      DOPBDOP : OUT std_logic_vector (1 DOWNTO 0) ;
      ADDRAWRADDR : IN std_logic_vector (12 DOWNTO 0) ;
      ADDRBRDADDR : IN std_logic_vector (12 DOWNTO 0) ;
      CLKAWRCLK : IN std_logic ;
      CLKBRDCLK : IN std_logic ;
      DIADI : IN std_logic_vector (15 DOWNTO 0) ;
      DIBDI : IN std_logic_vector (15 DOWNTO 0) ;
      DIPADIP : IN std_logic_vector (1 DOWNTO 0) ;
      DIPBDIP : IN std_logic_vector (1 DOWNTO 0) ;
      ENAWREN : IN std_logic ;
      ENBRDEN : IN std_logic ;
      REGCEA : IN std_logic ;
      REGCEBREGCE : IN std_logic ;
      RSTA : IN std_logic ;
      RSTBRST : IN std_logic ;
      WEAWEL : IN std_logic_vector (1 DOWNTO 0) ;
      WEBWEU : IN std_logic_vector (1 DOWNTO 0)) ;
   attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      RAMB8BWER : entity is true;
      end RAMB8BWER ;

architecture NETLIST of RAMB8BWER is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  RAMB16BWER
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity RAMB16BWER is 
   generic (DATA_WIDTH_A : integer := 0;
      DATA_WIDTH_B : integer := 0;
      DOA_REG : integer := 0;
      DOB_REG : integer := 0;
      EN_RSTRAM_A : boolean := TRUE;
      EN_RSTRAM_B : boolean := TRUE
      ;
      INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
      ;
      INIT_A : bit_vector := X"000000000"
      ;
      INIT_B : bit_vector := X"000000000";
      INIT_FILE : string := "NONE";
      RSTTYPE : string := "SYNC";
      RST_PRIORITY_A : string := "CE";
      RST_PRIORITY_B : string := "CE";
      SETUP_ALL : time := 1000000 ns;
      SETUP_READ_FIRST : time := 3000000 ns
      ;
      SIM_COLLISION_CHECK : string := "ALL"
      ;
      SIM_DEVICE : string := "SPARTAN3ADSP"
      ;
      SRVAL_A : bit_vector := X"000000000"
      ;
      SRVAL_B : bit_vector := X"000000000"
      ;
      WRITE_MODE_A : string := "WRITE_FIRST"
      ;
      WRITE_MODE_B : string := "WRITE_FIRST") ;
   
   port (
      DOA : OUT std_logic_vector (31 DOWNTO 0) ;
      DOB : OUT std_logic_vector (31 DOWNTO 0) ;
      DOPA : OUT std_logic_vector (3 DOWNTO 0) ;
      DOPB : OUT std_logic_vector (3 DOWNTO 0) ;
      ADDRA : IN std_logic_vector (13 DOWNTO 0) ;
      ADDRB : IN std_logic_vector (13 DOWNTO 0) ;
      CLKA : IN std_logic ;
      CLKB : IN std_logic ;
      DIA : IN std_logic_vector (31 DOWNTO 0) ;
      DIB : IN std_logic_vector (31 DOWNTO 0) ;
      DIPA : IN std_logic_vector (3 DOWNTO 0) ;
      DIPB : IN std_logic_vector (3 DOWNTO 0) ;
      ENA : IN std_logic ;
      ENB : IN std_logic ;
      REGCEA : IN std_logic ;
      REGCEB : IN std_logic ;
      RSTA : IN std_logic ;
      RSTB : IN std_logic ;
      WEA : IN std_logic_vector (3 DOWNTO 0) ;
      WEB : IN std_logic_vector (3 DOWNTO 0)) ;
   attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      RAMB16BWER : entity is true;
      end RAMB16BWER ;

architecture NETLIST of RAMB16BWER is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  FIFO18
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity FIFO18 is 
   generic (ALMOST_EMPTY_OFFSET : bit_vector := X"080"
      ;
      ALMOST_FULL_OFFSET : bit_vector := X"080";
      DATA_WIDTH : integer := 4;
      DO_REG : integer := 1;
      EN_SYN : boolean := FALSE;
      FIRST_WORD_FALL_THROUGH : boolean := FALSE
      ;
      SIM_MODE : string := "SAFE") ;
   
   port (
      ALMOSTEMPTY : OUT std_logic ;
      ALMOSTFULL : OUT std_logic ;
      DO : OUT std_logic_vector (15 DOWNTO 0) ;
      DOP : OUT std_logic_vector (1 DOWNTO 0) ;
      EMPTY : OUT std_logic ;
      FULL : OUT std_logic ;
      RDCOUNT : OUT std_logic_vector (11 DOWNTO 0) ;
      RDERR : OUT std_logic ;
      WRCOUNT : OUT std_logic_vector (11 DOWNTO 0) ;
      WRERR : OUT std_logic ;
      DI : IN std_logic_vector (15 DOWNTO 0) ;
      DIP : IN std_logic_vector (1 DOWNTO 0) ;
      RDCLK : IN std_logic ;
      RDEN : IN std_logic ;
      RST : IN std_logic ;
      WRCLK : IN std_logic ;
      WREN : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      FIFO18 : entity is true;
      end FIFO18 ;

architecture NETLIST of FIFO18 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  FIFO18_36
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity FIFO18_36 is 
   generic (ALMOST_EMPTY_OFFSET : bit_vector := X"080"
      ;
      ALMOST_FULL_OFFSET : bit_vector := X"080";
      DO_REG : integer := 1;
      EN_SYN : boolean := FALSE;
      FIRST_WORD_FALL_THROUGH : boolean := FALSE
      ;
      SIM_MODE : string := "SAFE") ;
   
   port (
      ALMOSTEMPTY : OUT std_logic ;
      ALMOSTFULL : OUT std_logic ;
      DO : OUT std_logic_vector (31 DOWNTO 0) ;
      DOP : OUT std_logic_vector (3 DOWNTO 0) ;
      EMPTY : OUT std_logic ;
      FULL : OUT std_logic ;
      RDCOUNT : OUT std_logic_vector (8 DOWNTO 0) ;
      RDERR : OUT std_logic ;
      WRCOUNT : OUT std_logic_vector (8 DOWNTO 0) ;
      WRERR : OUT std_logic ;
      DI : IN std_logic_vector (31 DOWNTO 0) ;
      DIP : IN std_logic_vector (3 DOWNTO 0) ;
      RDCLK : IN std_logic ;
      RDEN : IN std_logic ;
      RST : IN std_logic ;
      WRCLK : IN std_logic ;
      WREN : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      FIFO18_36 : entity is true;
      end FIFO18_36 ;

architecture NETLIST of FIFO18_36 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  FIFO36
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity FIFO36 is 
   generic (ALMOST_EMPTY_OFFSET : bit_vector := X"0080"
      ;
      ALMOST_FULL_OFFSET : bit_vector := X"0080";
      DATA_WIDTH : integer := 4;
      DO_REG : integer := 1;
      EN_SYN : boolean := FALSE;
      FIRST_WORD_FALL_THROUGH : boolean := FALSE
      ;
      SIM_MODE : string := "SAFE") ;
   
   port (
      ALMOSTEMPTY : OUT std_logic ;
      ALMOSTFULL : OUT std_logic ;
      DO : OUT std_logic_vector (31 DOWNTO 0) ;
      DOP : OUT std_logic_vector (3 DOWNTO 0) ;
      EMPTY : OUT std_logic ;
      FULL : OUT std_logic ;
      RDCOUNT : OUT std_logic_vector (12 DOWNTO 0) ;
      RDERR : OUT std_logic ;
      WRCOUNT : OUT std_logic_vector (12 DOWNTO 0) ;
      WRERR : OUT std_logic ;
      DI : IN std_logic_vector (31 DOWNTO 0) ;
      DIP : IN std_logic_vector (3 DOWNTO 0) ;
      RDCLK : IN std_logic ;
      RDEN : IN std_logic ;
      RST : IN std_logic ;
      WRCLK : IN std_logic ;
      WREN : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      FIFO36 : entity is true;
      end FIFO36 ;

architecture NETLIST of FIFO36 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  FIFO36_72
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity FIFO36_72 is 
   generic (ALMOST_EMPTY_OFFSET : bit_vector := X"080"
      ;
      ALMOST_FULL_OFFSET : bit_vector := X"080";
      DO_REG : integer := 1;
      EN_ECC_READ : boolean := FALSE;
      EN_ECC_WRITE : boolean := FALSE;
      EN_SYN : boolean := FALSE;
      FIRST_WORD_FALL_THROUGH : boolean := FALSE
      ;
      SIM_MODE : string := "SAFE") ;
   
   port (
      ALMOSTEMPTY : OUT std_logic ;
      ALMOSTFULL : OUT std_logic ;
      DBITERR : OUT std_logic ;
      DO : OUT std_logic_vector (63 DOWNTO 0) ;
      DOP : OUT std_logic_vector (7 DOWNTO 0) ;
      ECCPARITY : OUT std_logic_vector (7 DOWNTO 0) ;
      EMPTY : OUT std_logic ;
      FULL : OUT std_logic ;
      RDCOUNT : OUT std_logic_vector (8 DOWNTO 0) ;
      RDERR : OUT std_logic ;
      SBITERR : OUT std_logic ;
      WRCOUNT : OUT std_logic_vector (8 DOWNTO 0) ;
      WRERR : OUT std_logic ;
      DI : IN std_logic_vector (63 DOWNTO 0) ;
      DIP : IN std_logic_vector (7 DOWNTO 0) ;
      RDCLK : IN std_logic ;
      RDEN : IN std_logic ;
      RST : IN std_logic ;
      WRCLK : IN std_logic ;
      WREN : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      FIFO36_72 : entity is true;
      end FIFO36_72 ;

architecture NETLIST of FIFO36_72 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  FIFO18E1
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity FIFO18E1 is 
   generic (ALMOST_EMPTY_OFFSET : bit_vector := X"0080"
      ;
      ALMOST_FULL_OFFSET : bit_vector := X"0080";
      DATA_WIDTH : integer := 4;
      DO_REG : integer := 1;
      EN_SYN : boolean := FALSE;
      FIFO_MODE : string := "FIFO18"
      ;
      FIRST_WORD_FALL_THROUGH : boolean := FALSE
      ;
      INIT : bit_vector := X"000000000";
      SIM_DEVICE : string := "VIRTEX6";
      SRVAL : bit_vector := X"000000000") ;
   
   port (
      ALMOSTEMPTY : OUT std_logic ;
      ALMOSTFULL : OUT std_logic ;
      DO : OUT std_logic_vector (31 DOWNTO 0) ;
      DOP : OUT std_logic_vector (3 DOWNTO 0) ;
      EMPTY : OUT std_logic ;
      FULL : OUT std_logic ;
      RDCOUNT : OUT std_logic_vector (11 DOWNTO 0) ;
      RDERR : OUT std_logic ;
      WRCOUNT : OUT std_logic_vector (11 DOWNTO 0) ;
      WRERR : OUT std_logic ;
      DI : IN std_logic_vector (31 DOWNTO 0) ;
      DIP : IN std_logic_vector (3 DOWNTO 0) ;
      RDCLK : IN std_logic ;
      RDEN : IN std_logic ;
      REGCE : IN std_logic ;
      RST : IN std_logic ;
      RSTREG : IN std_logic ;
      WRCLK : IN std_logic ;
      WREN : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      FIFO18E1 : entity is true;
      end FIFO18E1 ;

architecture NETLIST of FIFO18E1 is       
      begin
      end NETLIST ;
      

-- 
-- Definition of  FIFO36E1
-- 
--      05/06/20 13:04:23
--      
--      Precision RTL Synthesis, 64-bit 2017.2.0.12
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Timing.all;

entity FIFO36E1 is 
   generic (ALMOST_EMPTY_OFFSET : BIT_VECTOR := X"0000010000000"
      ;
      ALMOST_FULL_OFFSET : BIT_VECTOR := X"0000010000000"
      ;
      DATA_WIDTH : INTEGER := 4;
      DO_REG : INTEGER := 1;
      EN_ECC_READ : STRING := "FALSE";
      EN_ECC_WRITE : STRING := "FALSE";
      EN_SYN : STRING := "FALSE";
      FIFO_MODE : STRING := "FIFO36"
      ;
      FIRST_WORD_FALL_THROUGH : STRING := "FALSE"
      ;
      INIT : BIT_VECTOR := X"000000000000000000000000000000000000000000000000000000000000000000000000"
      ;
      IS_RDCLK_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_RDEN_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_RSTREG_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_RST_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_WRCLK_INVERTED : BIT_VECTOR := X"0"
      ;
      IS_WREN_INVERTED : BIT_VECTOR := X"0"
      ;
      SIM_DEVICE : STRING := "7SERIES"
      ;
      SRVAL : BIT_VECTOR := X"000000000000000000000000000000000000000000000000000000000000000000000000"
   ) ;
   
   port (
      ALMOSTEMPTY : OUT std_logic ;
      ALMOSTFULL : OUT std_logic ;
      DBITERR : OUT std_logic ;
      DO : OUT std_logic_vector (63 DOWNTO 0) ;
      DOP : OUT std_logic_vector (7 DOWNTO 0) ;
      ECCPARITY : OUT std_logic_vector (7 DOWNTO 0) ;
      EMPTY : OUT std_logic ;
      FULL : OUT std_logic ;
      RDCOUNT : OUT std_logic_vector (12 DOWNTO 0) ;
      RDERR : OUT std_logic ;
      SBITERR : OUT std_logic ;
      WRCOUNT : OUT std_logic_vector (12 DOWNTO 0) ;
      WRERR : OUT std_logic ;
      DI : IN std_logic_vector (63 DOWNTO 0) ;
      DIP : IN std_logic_vector (7 DOWNTO 0) ;
      INJECTDBITERR : IN std_logic ;
      INJECTSBITERR : IN std_logic ;
      RDCLK : IN std_logic ;
      RDEN : IN std_logic ;
      REGCE : IN std_logic ;
      RST : IN std_logic ;
      RSTREG : IN std_logic ;
      WRCLK : IN std_logic ;
      WREN : IN std_logic) ;attribute RTLC_TECH_CELL: boolean;
   attribute RTLC_TECH_CELL of 
      FIFO36E1 : entity is true;
      end FIFO36E1 ;

architecture NETLIST of FIFO36E1 is       
      begin
      end NETLIST ;
      
