//
// Verilog Module Ethernet.V1
//
// Created:
//          by - waly.UNKNOWN (EGC-WALY-LT)
//          at - 02:40:29 05/13/2020
//
// using Mentor Graphics HDL Designer(TM) 2020.2 Built on 2 Mar 2020 at 18:07:13
//

`resetall
`timescale 1ns/10ps
module V1 ;


// ### Please start your Verilog code here ### 

endmodule
